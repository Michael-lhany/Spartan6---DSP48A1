module DSP_tb ();
reg CEA,CEB,CEC,CED,CEM,CEOPMODE,CEP,RSTA,RSTB,RSTC,RSTD,RSTM,RSTOPMODE,RSTP,RSTCARRYIN,CARRYIN,CLK,CECARRYIN;
reg [17:0] A,B,D,BCIN;
reg [47:0] C,PCIN;
reg [7:0] OPMODE;
wire CARRYOUT,CARRYOUTF;
wire [17:0] BCOUT;
wire [35:0] M;
wire [47:0] P, PCOUT;
parameter A0REG=0, A1REG=1, B0REG=0, B1REG=1, CREG=1, DREG=1,
		  MREG=1, PREG=1, CARRYINREG=1, CARRYOUTREG=1, OPMODEREG=1,
		  CARRYINSEL="OPMODE5",B_INPUT="DIRECT",RSSTYPE="SYNC";
DSP #(.A0REG(A0REG),.A1REG(A1REG),.B0REG(B0REG),.B1REG(B1REG),.CREG(CREG),.DREG(DREG),.MREG(MREG),.PREG(PREG),.CARRYINREG(CARRYINREG),
	.CARRYOUTREG(CARRYOUTREG),.OPMODEREG(OPMODEREG),.CARRYINSEL(CARRYINSEL),.B_INPUT(B_INPUT),.RSSTYPE(RSSTYPE)) dut (A,B,C,D,CARRYIN,
	M,P,CARRYOUT,CARRYOUTF,CLK,OPMODE,CEA,CEB,CEC,CED,CEM,CEOPMODE,CECARRYIN,CEP,RSTA,RSTB,RSTC,RSTD,RSTM,RSTOPMODE,RSTP,RSTCARRYIN,BCIN,BCOUT,PCIN,PCOUT);
initial		begin
	CLK=0;
	forever
	#1	CLK=~CLK;
end
integer i;
initial begin
	CEA=1;
	CEB=1;
	CEC=1;
	CED=1;
	CEM=1;
	CEOPMODE=1;
	CEP=1;
	RSTA=0;RSTB=0;RSTC=0;RSTD=0;RSTM=0;RSTOPMODE=0;RSTP=0;
	RSTCARRYIN=0;CECARRYIN=1;
	for (i = 0; i < 20; i=i+1) begin
		OPMODE=$random;
		CARRYIN=$random;A=$random;B=$random;
		D=$random;BCIN=$random;C=$random;
		PCIN=$random;
		#8;
	end
	$stop;
end
endmodule